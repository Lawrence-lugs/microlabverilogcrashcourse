module ALU (
    input [3:0] a, b,
    input [2:0] opcode,
    output reg [3:0] result,
    output reg zero
);

    // TODO: Do your stuff!

endmodule