`timescale 1ns/1ps

module tb_queue;

// Write the testbench here

endmodule