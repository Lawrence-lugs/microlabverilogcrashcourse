`timescale 1ns/1ps

module tb_queue;

    // Write your testbench here

    // Make sure to test the following
    // 1. Enqueue and Dequeue operations
    // 2. Full and Empty conditions
    // 3. Enqueue when full, Dequeue when empty

endmodule